module job_q_2.8(
  input [3:0] A, 
  input [3:0] B, 
  output [3:0] Sum
);
  assign Sum = A + B;
endmodule
